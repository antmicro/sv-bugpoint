`verilator_config
// irremovable verilator_config section
