module full_adder (
        input cin);
endmodule
