module t;
endmodule