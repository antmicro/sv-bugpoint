module t;
    initial begin
        $finish;
    end
endmodule
