

module full_adder3 (
        input cin);
endmodule
