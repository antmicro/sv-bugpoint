package doe_defines_pkg;  
typedef enum logic [1:0] {
    DOE_NOP    = 2'b00
} doe_cmd_e;
endpackage
