module t;
  initial begin;
    $finish;
  end;
endmodule
// irremovable comment with no newline