// nonsense code that should error out on access to undefined struct member

module full_adder (
        input a,
        input b,
        input cin,
        output s,
        output cout);
    assign s = a^b^cin;
    assign cout = (a&b) | (b&cin) | (a&cin);
endmodule

module full_adder2 (
        input a,
        input b,
        input cin,
        output s,
        output cout);
    assign s = a^b^cin;
    assign cout = (a&b) | (b&cin) | (a&cin);
endmodule

module full_adder3 (
        input a,
        input b,
        input cin,
        output s,
        output cout);
    assign s = a^b^cin;
    assign cout = (a&b) | (b&cin) | (a&cin);
endmodule

typedef struct {
        byte a;
        int b;
} struct_foo;

module serial_adder #(WIDTH=32) (
        input  [WIDTH-1:0] a,
        input  [WIDTH-1:0] b,
        input  cin,
        output [WIDTH-1:0] s,
        output cout);

    wire [WIDTH:0] k;
    wire [WIDTH:0] l;
    wire [WIDTH:0] c;
    wire [WIDTH:0] m;
    wire [WIDTH:0] n = 4;

    generate for (genvar i = 0; i < WIDTH; i++)
        full_adder fa(a[i], b[i], c[i], s[i], c[i+1]);
    endgenerate


    struct_foo foo = '{5,6};
    assign foo.a = 25;

    wire [3:0] x = 4'hF;
    wire [3:0] y = 5'h1F;
    
    assign c[0] = cin;
    assign cout = c[WIDTH];

endmodule

