module t;
    initial begin: label
        $finish;
    end: label
endmodule : t
