../examples/caliptra_vcd/sv-bugpoint-input.sv