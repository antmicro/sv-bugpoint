// non-functional comment, should be removed
`verilator_config
// irremovable verilator_config section
