// irremovable comment with no newline